----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:24:14 05/19/2007 
-- Design Name: 
-- Module Name:    Comp8 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Comp24 is
    Port ( FN1 : in  STD_ULOGIC_VECTOR (23 downto 0);
           FN2 : in  STD_ULOGIC_VECTOR (23 downto 0);
           S, EQ : out  STD_ULOGIC);
end Comp24;

architecture Behavioral of Comp24 is
signal X:std_Ulogic_vector(23 downto 0);

begin

X(23)<= FN1(23) XNOR FN2(23);
X(22)<= FN1(22) XNOR FN2(22);
X(21)<= FN1(21) XNOR FN2(21);
X(20)<= FN1(20) XNOR FN2(20);
X(19)<= FN1(19) XNOR FN2(19);
X(18)<= FN1(18) XNOR FN2(18);
X(17)<= FN1(17) XNOR FN2(17);
X(16)<= FN1(16) XNOR FN2(16);
X(15)<= FN1(15) XNOR FN2(15);
X(14)<= FN1(14) XNOR FN2(14);
X(13)<= FN1(13) XNOR FN2(13);
X(12)<= FN1(12) XNOR FN2(12);
X(11)<= FN1(11) XNOR FN2(11);
X(10)<= FN1(10) XNOR FN2(10);
X(9)<= FN1(9) XNOR FN2(9);
X(8)<= FN1(8) XNOR FN2(8);
X(7)<= FN1(7) XNOR FN2(7);
X(6)<= FN1(6) XNOR FN2(6);
X(5)<= FN1(5) XNOR FN2(5);
X(4)<= FN1(4) XNOR FN2(4);
X(3)<= FN1(3) XNOR FN2(3);
X(2)<= FN1(2) XNOR FN2(2);
X(1)<= FN1(1) XNOR FN2(1);
X(0)<= FN1(0) XNOR FN2(0);

S <= ((NOT FN1(23)) AND FN2(23)) 
		OR (X(23)AND(NOT FN1(22)) AND FN2(22)) 
		OR (X(23)AND X(22)AND(NOT FN1(21)) AND FN2(21)) 
		OR (X(23)AND X(22)AND X(21)AND(NOT FN1(20)) AND FN2(20))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND(NOT FN1(19)) AND FN2(19)) 
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND(NOT FN1(18)) AND FN2(18))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND(NOT FN1(17)) AND FN2(17))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND(NOT FN1(16)) AND FN2(16))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND(NOT FN1(15)) AND FN2(15))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND(NOT FN1(14)) AND FN2(14))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND(NOT FN1(13)) AND FN2(13))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND X(13)AND(NOT FN1(12)) AND FN2(12))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND X(13)AND X(12)AND(NOT FN1(11)) AND FN2(11))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND X(13)AND X(12)AND X(11)AND(NOT FN1(10)) AND FN2(10))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND X(13)AND X(12)AND X(11)AND X(10)AND(NOT FN1(9)) AND FN2(9))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND X(13)AND X(12)AND X(11)AND X(10)AND X(9)AND(NOT FN1(8)) AND FN2(8))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND X(13)AND X(12)AND X(11)AND X(10)AND X(9)AND X(8)AND(NOT FN1(7)) AND FN2(7))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND X(13)AND X(12)AND X(11)AND X(10)AND X(9)AND X(8)AND X(7)AND(NOT FN1(6)) AND FN2(6))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND X(13)AND X(12)AND X(11)AND X(10)AND X(9)AND X(8)AND X(7)AND X(6)AND(NOT FN1(5)) AND FN2(5))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND X(13)AND X(12)AND X(11)AND X(10)AND X(9)AND X(8)AND X(7)AND X(6)AND X(5)AND(NOT FN1(4)) AND FN2(4))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND X(13)AND X(12)AND X(11)AND X(10)AND X(9)AND X(8)AND X(7)AND X(6)AND X(5)AND X(4)AND(NOT FN1(3)) AND FN2(3))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND X(13)AND X(12)AND X(11)AND X(10)AND X(9)AND X(8)AND X(7)AND X(6)AND X(5)AND X(4)AND X(3)AND(NOT FN1(2)) AND FN2(2))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND X(13)AND X(12)AND X(11)AND X(10)AND X(9)AND X(8)AND X(7)AND X(6)AND X(5)AND X(4)AND X(3)AND X(2)AND(NOT FN1(1)) AND FN2(1))
		OR (X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND X(13)AND X(12)AND X(11)AND X(10)AND X(9)AND X(8)AND X(7)AND X(6)AND X(5)AND X(4)AND X(3)AND X(2)AND X(1)AND(NOT FN1(0)) AND FN2(0));
		
		EQ <= X(23)AND X(22)AND X(21)AND X(20)AND X(19)AND X(18)AND X(17)AND X(16)AND X(15)AND X(14)AND X(13)AND X(12)AND X(11)AND X(10)AND X(9)AND X(8)AND X(7)AND X(6)AND X(5)AND X(4)AND X(3)AND X(2)AND X(1)AND X(0);
end Behavioral;
